// ------------------------------------------------------------------------- 
// File name    : AHB_UVC_checker_c.sv
// Title        : AHB_UVC Checker
// Project      : AHB_UVC 
// Created On   : 2024-02-07
// Developers   : 
// -------------------------------------------------------------------------

`ifndef AHB_UVC_CHECKER_SV
`define AHB_UVC_CHECKER_SV
interface AHB_UVC_checker;
endinterface : AHB_UVC_checker
`endif

